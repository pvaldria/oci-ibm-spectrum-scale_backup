ss-server-5.privateb0.gpfs.oraclevcn.com slots=52
ss-server-6.privateb0.gpfs.oraclevcn.com slots=52
